bind top_zynq license_guard u_license_enforcer();

